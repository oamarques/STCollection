    5
    1.0
    2.0
    3.0
    4.0
    5.0
