      20
   10.23838
   10.23838
    9.05117
    9.05117
    8.03258
    8.03258
    7.03589
    7.03589
    6.04188
    6.04188
    5.05037
    5.05037
    4.06324
    4.06322
    3.08626
    3.08397
    2.17808
    2.08889
    1.41732
    0.50883
