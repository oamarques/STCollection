    5
    1.5
    2.8
    2.8
    2.8
    4.6
