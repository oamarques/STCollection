    5
    1.5
    2.8
    0.0
    3.6
    4.6
