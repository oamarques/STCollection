      40
   20.23177
   20.23177
   19.03659
   19.03659
   18.01505
   18.01505
   17.01474
   17.01474
   16.01564
   16.01564
   15.01668
   15.01668
   14.01787
   14.01787
   13.01925
   13.01925
   12.02086
   12.02086
   11.02276
   11.02276
   10.02505
   10.02505
    9.02784
    9.02784
    8.03134
    8.03134
    7.03585
    7.03585
    6.04188
    6.04188
    5.05037
    5.05037
    4.06324
    4.06322
    3.08626
    3.08397
    2.17808
    2.08889
    1.41732
    0.50883
