      30
   15.23394
   15.23394
   14.04127
   14.04127
   13.02043
   13.02043
   12.02089
   12.02089
   11.02276
   11.02276
   10.02505
   10.02505
    9.02784
    9.02784
    8.03134
    8.03134
    7.03585
    7.03585
    6.04188
    6.04188
    5.05037
    5.05037
    4.06324
    4.06322
    3.08626
    3.08397
    2.17808
    2.08889
    1.41732
    0.50883
